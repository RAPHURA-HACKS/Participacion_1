//1.Definicion del modulo, sus entradas y salidas
//Dentro del parentesis se define los 1/0
module _and (input a, input b, output c);
//2.Definen cables o componentes internos
//N/A
//3.Asignaciones, instancias y conexiones

assign c= a & b;
endmodule